module InsMem (
    addr,
    datain,
    dataout,
    sigwr,
    sigon,
    clk
);
  input [6:0] addr;
  input [31:0] datain;
  output reg [31:0] dataout;
  input sigwr;
  input sigon;
  input clk;

  reg [31:0] mem[127:0];

  initial begin
    mem[0]  <= 32'b00000100001000000000000000011000;
    mem[1]  <= 32'b01001100000000010000000000000000;
    mem[2]  <= 32'b01111000000000010000000000000000;
    mem[3]  <= 32'b00000100001000000000000000101101;
    mem[4]  <= 32'b01001100000000010000000000000001;
    mem[5]  <= 32'b01111000000000010000000000000000;
    mem[6]  <= 32'b00000100001000000000000000001010;
    mem[7]  <= 32'b01001100000000010000000000000010;
    mem[8]  <= 32'b01111000000000010000000000000000;
    mem[9]  <= 32'b00000100001000000000000000001000;
    mem[10] <= 32'b01001100000000010000000000000011;
    mem[11] <= 32'b01111000000000010000000000000000;
    mem[12] <= 32'b00000100001000000000000000010110;
    mem[13] <= 32'b01001100000000010000000000000100;
    mem[14] <= 32'b01111000000000010000000000000000;
    mem[15] <= 32'b00000100001111111111111110011100;
    mem[16] <= 32'b01001100000000010000000000000101;
    mem[17] <= 32'b01111000000000010000000000000000;
    mem[18] <= 32'b00000100001111111111111111011110;
    mem[19] <= 32'b01001100000000010000000000000110;
    mem[20] <= 32'b01111000000000010000000000000000;
    mem[21] <= 32'b00000100001000000000000001011010;
    mem[22] <= 32'b01001100000000010000000000000111;
    mem[23] <= 32'b01111000000000010000000000000000;
    mem[24] <= 32'b00000100001000000000000000000000;
    mem[25] <= 32'b01001100000000010000000000001000;
    mem[26] <= 32'b01111000000000010000000000000000;
    mem[27] <= 32'b00000100001111111111111111101001;
    mem[28] <= 32'b01001100000000010000000000001001;
    mem[29] <= 32'b01111000000000010000000000000000;
    mem[30] <= 32'b00000100001000000000000000001000;
    mem[31] <= 32'b00000100010000000000000000001001;
    mem[32] <= 32'b00001100010000000000000000000001;
    mem[33] <= 32'b01011100010000000000000000010011;
    mem[34] <= 32'b00001000001000100001100000000000;
    mem[35] <= 32'b00001000001000110010000000000000;
    mem[36] <= 32'b01111000100001010000000000000000;
    mem[37] <= 32'b00000100101000000000000000000001;
    mem[38] <= 32'b00001100101000000000000000000001;
    mem[39] <= 32'b01011100101000000000000000001100;
    mem[40] <= 32'b00001000100001010011000000000000;
    mem[41] <= 32'b01001000110001110000000000000000;
    mem[42] <= 32'b01001000110010000000000000000001;
    mem[43] <= 32'b00001001000001110100100000000000;
    mem[44] <= 32'b01100001001000000000000000000110;
    mem[45] <= 32'b00000001000001110100000000000000;
    mem[46] <= 32'b00001001000001110011100000000000;
    mem[47] <= 32'b00001001000001110100000000000000;
    mem[48] <= 32'b01001100110001110000000000000000;
    mem[49] <= 32'b01001100110010000000000000000001;
    mem[50] <= 32'b01011011111111111111111111110100;
    mem[51] <= 32'b01011011111111111111111111101101;
  end

  always @(addr or datain or sigwr or sigon) begin
    if (sigon) begin
      if (sigwr) begin
        mem[addr] = datain;
        dataout   = datain;
      end else begin
        dataout = mem[addr];
      end
    end
  end
endmodule